LIBRARY ieee;
USE ieee.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;

--  Entity Declaration

ENTITY UartToRS IS
    -- {{ALTERA_IO_BEGIN}} DO NOT REMOVE THIS LINE!
    PORT
    (
    -------------------------------������������ ������-----------------------------------
        clk     :   in STD_LOGIC;                           -- 80.000.000 Hz
--------------------------------��Ȩ���� ������-------------------------------------
        RS485_RX        : in std_logic;                     -- �����
        data_out: out std_logic_vector (7 downto 0);        -- ����������
        RX_VALID: out std_logic                          -- �������
---------------------------------��Ȩ������������------------------------------------
        --inDreq  : in STD_LOGIC;                             -- ������ ������ ������� �� �����
       -- reqBus: in STD_LOGIC_VECTOR (0 to 9);             -- ��������� ����
       -- RS485_TX: out STD_LOGIC;                            -- ���������������� ������ �����������
        --dir_TX  : out STD_LOGIC;                            -- ������� �����������
        --dir_RX  : out STD_LOGIC;                             -- ����� � �������� ��������������
        --cnt_ram : out integer range 0 to 880
    );
    -- {{ALTERA_IO_END}} DO NOT REMOVE THIS LINE!
    
END UartToRS;


--  Architecture Body

ARCHITECTURE UartToRS_architecture OF UartToRS IS

signal rx_act   : std_logic;                                -- ��������������� ������ ���������� �����

signal clk5MHz  : STD_LOGIC;                                -- ���������� ������� 5 ��� ��� ������������ RS-485
signal TXenable : STD_LOGIC;                                -- ��������������� ������ ���������� ��������

BEGIN
process (clk, clk5MHz)
----------------------------------------------
----- ���������� ��� ��Ȩ����� �� UART  ------
----------------------------------------------
variable place  : integer range 0 to 8 := 0;                -- ����� ���� ���������� � ����������
variable data   : std_logic_vector (7 downto 0);            -- ���������� � �������
variable strtcnt: integer range 0 to 8 := 0;                -- ������� ���������� ����
variable stepcnt: integer range 0 to 16 := 0;               -- ������� ������ ����� ������
variable newcnt : integer range 0 to 10 := 0;
variable VALID	: std_logic;
----------------------------------------------

-----------------------------------------------------------------------------------------------------------------
-----------------------------------------------------------------------------------------------------------------
-----------------------------------------------------------------------------------------------------------------
begin
--RX_VALID <= VALID;                                                    --
----------------------------------------------
----- ������ ��Ȩ�����. ����� ����������  ----
----------------------------------------------
if rising_edge(clk) then
RX_VALID <= VALID; 
--    RX_VALID <= '0';                                        -- �������� �� ��������� ��������� ������������
	if(VALID = '1') then
		newcnt := newcnt + 1;
		if(newcnt = 10) then
			VALID := '0';
			newcnt := 0;
		end if;
	end if;
    if (RS485_RX = '0') and (rx_act = '0') then                 -- ����� ��������� ���
		
        strtcnt := strtcnt + 1;                             -- ��������� �������� ���������� ����
        --strcnt==4 ��� 40 ���
        if (strtcnt = 4) then                               --
            rx_act <= '1';                                  -- ����� ������� �������� ��������
            strtcnt := 0;                                   -- � ������� ������� ��� ��������� ��������
        end if;                                             --
    end if;
    if (rx_act = '1') then                                  -- ���� �������� ��������� ��������
        stepcnt := stepcnt + 1;                             -- ����� ������� ����� ��� ������� ����
         --stepcnt==8 ��� 40 ���
        if (stepcnt = 8)then                               -- �������� ����������
            if (place = 8) then                             -- � ����� �����, ���� ����� �� ������� ����������
                if (RS485_RX = '1') then                    -- ���� ����� ����-���
                    rx_act <= '0';                          -- ����� ������� �������� �����������
                    VALID := '1';                        -- ����� ������� �������� ����������
                    data_out <= data;                       -- �������� �� ���� ��������� ����������
                    place := 0;                             -- ������� ��������
                    stepcnt := 0;                           -- ���������� � ������
                else                                        -- � ��������� ������
                    rx_act <= '0';                          -- �������� ��������
                    place := 0;                             -- ������� ��������
                    stepcnt := 0;                           -- � �� ������ ����������
                end if;                                     -- ������� �������� �����
            else                                            -- � ���� � ��� �� ����� ��������, ��
                data(place) := RS485_RX;                    -- ������� � ���������� ������ �� �����
                place := place + 1;                         -- �������������� ����� � ����������
                stepcnt := 0;                               -- ������� ������� ������
            end if;                                         -- ��������� � ��� �� ����
        end if;                                             --
    end if;
end if;

end process;
END UartToRS_architecture;