// megafunction wizard: %LPM_MUX%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: lpm_mux 

// ============================================================
// File Name: MUXmem.v
// Megafunction Name(s):
// 			lpm_mux
//
// Simulation Library Files(s):
// 			lpm
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 9.0 Build 184 04/29/2009 SP 1 SJ Web Edition
// ************************************************************


//Copyright (C) 1991-2009 Altera Corporation
//Your use of Altera Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Altera Program License 
//Subscription Agreement, Altera MegaCore Function License 
//Agreement, or other applicable license agreement, including, 
//without limitation, that your use is for the sole purpose of 
//programming logic devices manufactured by Altera and sold by 
//Altera or its authorized distributors.  Please refer to the 
//applicable agreement for further details.


// synopsys translate_off
`timescale 1 ps / 1 ps
// synopsys translate_on
module MUXmem (
	data0x,
	data1x,
	data2x,
	sel,
	result);

	input	[17:0]  data0x;
	input	[17:0]  data1x;
	input	[17:0]  data2x;
	input	[1:0]  sel;
	output	[17:0]  result;

	wire [17:0] sub_wire0;
	wire [17:0] sub_wire4 = data2x[17:0];
	wire [17:0] sub_wire3 = data0x[17:0];
	wire [17:0] result = sub_wire0[17:0];
	wire [17:0] sub_wire1 = data1x[17:0];
	wire [53:0] sub_wire2 = {sub_wire4, sub_wire1, sub_wire3};

	lpm_mux	lpm_mux_component (
				.sel (sel),
				.data (sub_wire2),
				.result (sub_wire0)
				// synopsys translate_off
				,
				.aclr (),
				.clken (),
				.clock ()
				// synopsys translate_on
				);
	defparam
		lpm_mux_component.lpm_size = 3,
		lpm_mux_component.lpm_type = "LPM_MUX",
		lpm_mux_component.lpm_width = 18,
		lpm_mux_component.lpm_widths = 2;


endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "FLEX10KE"
// Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
// Retrieval info: CONSTANT: LPM_SIZE NUMERIC "3"
// Retrieval info: CONSTANT: LPM_TYPE STRING "LPM_MUX"
// Retrieval info: CONSTANT: LPM_WIDTH NUMERIC "18"
// Retrieval info: CONSTANT: LPM_WIDTHS NUMERIC "2"
// Retrieval info: USED_PORT: data0x 0 0 18 0 INPUT NODEFVAL data0x[17..0]
// Retrieval info: USED_PORT: data1x 0 0 18 0 INPUT NODEFVAL data1x[17..0]
// Retrieval info: USED_PORT: data2x 0 0 18 0 INPUT NODEFVAL data2x[17..0]
// Retrieval info: USED_PORT: result 0 0 18 0 OUTPUT NODEFVAL result[17..0]
// Retrieval info: USED_PORT: sel 0 0 2 0 INPUT NODEFVAL sel[1..0]
// Retrieval info: CONNECT: result 0 0 18 0 @result 0 0 18 0
// Retrieval info: CONNECT: @data 0 0 18 36 data2x 0 0 18 0
// Retrieval info: CONNECT: @data 0 0 18 18 data1x 0 0 18 0
// Retrieval info: CONNECT: @data 0 0 18 0 data0x 0 0 18 0
// Retrieval info: CONNECT: @sel 0 0 2 0 sel 0 0 2 0
// Retrieval info: LIBRARY: lpm lpm.lpm_components.all
// Retrieval info: GEN_FILE: TYPE_NORMAL MUXmem.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL MUXmem.inc FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL MUXmem.cmp TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL MUXmem.bsf TRUE FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL MUXmem_inst.v FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL MUXmem_bb.v TRUE
// Retrieval info: LIB_FILE: lpm
